module vacio();

endmodule 