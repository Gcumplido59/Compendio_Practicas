module topLevelSum(
	input x, y,
	output a,b,c,d,e,f,g,
	wire w0,w1;
);

adder u1();

decdisp u2();

endmodule